module MIPS_Pipeline_Top (
    input clk,
    input reset
);

    // ==============================================================================
    // CABLES (WIRES) DE INTERCONEXIÓN ENTRE ETAPAS
    // ==============================================================================

    // --- Etapa IF (Instruction Fetch) ---
    wire [31:0] pc_in, pc_out, pc_plus_4;
    wire [31:0] instr;
    wire [31:0] branch_target_address;
    wire pcsrc; // Selector para salto (Branch)

    // --- Etapa ID (Instruction Decode) ---
    wire [31:0] if_id_pc_next, if_id_instr;
    wire [31:0] read_data1, read_data2, sign_ext_imm;
    wire [4:0]  rs_addr, rt_addr, rd_addr;
    
    // Señales de Control puras (salida de la Control Unit)
    wire ctrl_reg_dst, ctrl_branch, ctrl_mem_read, ctrl_mem_to_reg;
    wire [1:0] ctrl_alu_op;
    wire ctrl_mem_write, ctrl_alu_src, ctrl_reg_write;
    
    // Cables para el Branch en ID (si pasamos el branch por buffers)
    wire id_ex_branch, ex_mem_branch;

    // --- Etapa EX (Execute) ---
    // Señales que salen del buffer ID/EX
    wire id_ex_reg_write, id_ex_mem_to_reg, id_ex_mem_read, id_ex_mem_write;
    wire id_ex_reg_dst, id_ex_alu_src;
    wire [1:0] id_ex_alu_op;
    wire [31:0] id_ex_pc_next, id_ex_read_data1, id_ex_read_data2, id_ex_sign_ext;
    wire [4:0]  id_ex_rs, id_ex_rt, id_ex_rd;
    
    // Cables internos de EX
    wire [31:0] alu_in_a, alu_in_b_temp, alu_in_b_final;
    wire [31:0] alu_result;
    wire zero_flag;
    wire [4:0]  write_reg_addr_ex; 
    wire [3:0]  alu_control_signal;
    wire [1:0]  forward_a, forward_b; // Del Forwarding Unit

    // --- Etapa MEM (Memory) ---
    // Señales que salen del buffer EX/MEM
    wire ex_mem_reg_write, ex_mem_mem_to_reg, ex_mem_mem_read, ex_mem_mem_write;
    wire ex_mem_zero; // Flag Zero viajando
    wire [31:0] ex_mem_alu_result, ex_mem_write_data;
    wire [4:0]  ex_mem_write_reg;
    wire [31:0] mem_read_data;

    // --- Etapa WB (Write Back) ---
    // Señales que salen del buffer MEM/WB
    wire mem_wb_reg_write, mem_wb_mem_to_reg;
    wire [31:0] mem_wb_read_data, mem_wb_alu_result;
    wire [4:0]  mem_wb_write_reg;
    wire [31:0] result_to_write; 

    // ==============================================================================
    // ETAPA 1: INSTRUCTION FETCH (IF)
    // ==============================================================================

    // Lógica básica de Branch: Si en la etapa MEM decidimos saltar
    assign pcsrc = ex_mem_branch & ex_mem_zero; 
    
    // Mux del PC (Branch vs PC+4)
    // NOTA: 'branch_target_address' debería calcularse correctamente. 
    // En este ejemplo simple asumimos que se calculó antes o se pasa el offset.
    // Para simplificar, aquí usaremos pc_plus_4 por defecto si no hay lógica de cálculo de branch completa.
    assign pc_in = (pcsrc) ? branch_target_address : pc_plus_4; 

    ProgramCounter PC (
        .clk(clk), .reset(reset), 
        .enable(1'b1), // SIEMPRE HABILITADO (Sin Hazard Unit)
        .pc_in(pc_in), .pc_out(pc_out)
    );

    Adder Add_PC4 (.a(pc_out), .b(32'd4), .result(pc_plus_4));

    InstructionMemory InstrMem (.address(pc_out), .instruction(instr));

    // ==============================================================================
    // BUFFER IF/ID
    // ==============================================================================
    IF_ID_Buffer IF_ID (
        .clk(clk), .reset(reset), 
        .enable(1'b1), // SIEMPRE HABILITADO (Sin Hazard Unit)
        .pc_next_in(pc_plus_4), .instr_in(instr),
        .pc_next_out(if_id_pc_next), .instr_out(if_id_instr)
    );

    // ==============================================================================
    // ETAPA 2: INSTRUCTION DECODE (ID)
    // ==============================================================================

    // >>> HAZARD UNIT ELIMINADA AQUÍ <<<

    ControlUnit Control (
        .opcode(if_id_instr[31:26]),
        .reg_dst(ctrl_reg_dst), .branch(ctrl_branch), .mem_read(ctrl_mem_read),
        .mem_to_reg(ctrl_mem_to_reg), .alu_op(ctrl_alu_op), .mem_write(ctrl_mem_write),
        .alu_src(ctrl_alu_src), .reg_write(ctrl_reg_write)
    );

    RegisterFile RegFile (
        .clk(clk), .reg_write(mem_wb_reg_write),
        .read_reg1(if_id_instr[25:21]), .read_reg2(if_id_instr[20:16]),
        .write_reg(mem_wb_write_reg), .write_data(result_to_write),
        .read_data1(read_data1), .read_data2(read_data2)
    );

    SignExtend SignExt (.in(if_id_instr[15:0]), .out(sign_ext_imm));

    // ==============================================================================
    // BUFFER ID/EX
    // ==============================================================================
    ID_EX_Buffer ID_EX (
        .clk(clk), .reset(reset),
        // Control (Directo, sin MUX de Hazard)
        .RegWrite_in(ctrl_reg_write),
        .MemtoReg_in(ctrl_mem_to_reg),
        .MemRead_in(ctrl_mem_read),
        .MemWrite_in(ctrl_mem_write),
        .RegDst_in(ctrl_reg_dst),
        .ALUSrc_in(ctrl_alu_src),
        .ALUOp_in(ctrl_alu_op),
        .Branch_in(ctrl_branch), // Conectado directo
        
        // Datos
        .pc_next_in(if_id_pc_next), .read_data1_in(read_data1), .read_data2_in(read_data2),
        .sign_ext_in(sign_ext_imm),
        .rs_in(if_id_instr[25:21]), .rt_in(if_id_instr[20:16]), .rd_in(if_id_instr[15:11]),
        
        // Salidas
        .RegWrite_out(id_ex_reg_write), .MemtoReg_out(id_ex_mem_to_reg),
        .MemRead_out(id_ex_mem_read), .MemWrite_out(id_ex_mem_write),
        .RegDst_out(id_ex_reg_dst), .ALUSrc_out(id_ex_alu_src), .ALUOp_out(id_ex_alu_op),
        .Branch_out(id_ex_branch),
        
        .pc_next_out(id_ex_pc_next), .read_data1_out(id_ex_read_data1), .read_data2_out(id_ex_read_data2),
        .sign_ext_out(id_ex_sign_ext),
        .rs_out(id_ex_rs), .rt_out(id_ex_rt), .rd_out(id_ex_rd)
    );

    // ==============================================================================
    // ETAPA 3: EXECUTE (EX)
    // ==============================================================================

    // Forwarding Unit (Se mantiene para dependencias de datos básicas)
    ForwardingUnit Forwarding (
        .ID_EX_Rs(id_ex_rs), .ID_EX_Rt(id_ex_rt),
        .EX_MEM_Rd(ex_mem_write_reg), .EX_MEM_RegWrite(ex_mem_reg_write),
        .MEM_WB_Rd(mem_wb_write_reg), .MEM_WB_RegWrite(mem_wb_reg_write),
        .ForwardA(forward_a), .ForwardB(forward_b)
    );

    // Muxes de Forwarding
    assign alu_in_a = (forward_a == 2'b10) ? ex_mem_alu_result :
                      (forward_a == 2'b01) ? result_to_write : id_ex_read_data1;

    assign alu_in_b_temp = (forward_b == 2'b10) ? ex_mem_alu_result :
                           (forward_b == 2'b01) ? result_to_write : id_ex_read_data2;

    assign alu_in_b_final = (id_ex_alu_src) ? id_ex_sign_ext : alu_in_b_temp;

    assign write_reg_addr_ex = (id_ex_reg_dst) ? id_ex_rd : id_ex_rt;

    // Cálculo de dirección de Branch (Shift + Add)
    // Nota: Necesitas instanciar aquí tu ShiftLeft2 y Adder si quieres calcular el salto
    // assign branch_target_address = id_ex_pc_next + (id_ex_sign_ext << 2); 
    // Por simplicidad lo dejo como wire, asegúrate de conectarlo si usas branches.

    ALUControl ALU_Ctrl (.alu_op(id_ex_alu_op), .funct(id_ex_sign_ext[5:0]), .alu_control_out(alu_control_signal));

    ALU Main_ALU (
        .a(alu_in_a), .b(alu_in_b_final), .alu_control(alu_control_signal),
        .result(alu_result), .zero(zero_flag)
    );

    // ==============================================================================
    // BUFFER EX/MEM
    // ==============================================================================
    EX_MEM_Buffer EX_MEM (
        .clk(clk), .reset(reset),
        .RegWrite_in(id_ex_reg_write), .MemtoReg_in(id_ex_mem_to_reg),
        .MemRead_in(id_ex_mem_read), .MemWrite_in(id_ex_mem_write),
        .Branch_in(id_ex_branch),
        
        .alu_result_in(alu_result), .write_data_in(alu_in_b_temp), 
        .write_reg_in(write_reg_addr_ex),
        .Zero_in(zero_flag),
        
        // Salidas
        .RegWrite_out(ex_mem_reg_write), .MemtoReg_out(ex_mem_mem_to_reg),
        .MemRead_out(ex_mem_mem_read), .MemWrite_out(ex_mem_mem_write),
        .Branch_out(ex_mem_branch),
        .Zero_out(ex_mem_zero),
        
        .alu_result_out(ex_mem_alu_result), .write_data_out(ex_mem_write_data),
        .write_reg_out(ex_mem_write_reg)
    );

    // ==============================================================================
    // ETAPA 4: MEMORY (MEM)
    // ==============================================================================

    DataMemory DataMem (
        .clk(clk), .address(ex_mem_alu_result),
        .write_data(ex_mem_write_data),
        .mem_write(ex_mem_mem_write), .mem_read(ex_mem_mem_read),
        .read_data(mem_read_data)
    );

    // ==============================================================================
    // BUFFER MEM/WB
    // ==============================================================================
    MEM_WB_Buffer MEM_WB (
        .clk(clk), .reset(reset),
        .RegWrite_in(ex_mem_reg_write), .MemtoReg_in(ex_mem_mem_to_reg),
        .mem_read_data_in(mem_read_data), .alu_result_in(ex_mem_alu_result),
        .write_reg_in(ex_mem_write_reg),
        // Salidas
        .RegWrite_out(mem_wb_reg_write), .MemtoReg_out(mem_wb_mem_to_reg),
        .mem_read_data_out(mem_wb_read_data), .alu_result_out(mem_wb_alu_result),
        .write_reg_out(mem_wb_write_reg)
    );

    // ==============================================================================
    // ETAPA 5: WRITE BACK (WB)
    // ==============================================================================

    assign result_to_write = (mem_wb_mem_to_reg) ? mem_wb_read_data : mem_wb_alu_result;

endmodule